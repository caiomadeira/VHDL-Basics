--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity soma_sub4 is
	port (-- <COMPLETAR>
	     );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture soma_sub4 of soma_sub4 is
	-- <COMPLETAR>
begin

    -- <COMPLETAR>

end architecture;