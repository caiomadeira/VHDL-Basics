--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity soma_sub8 is
	port (-- <COMPLETAR>
	     );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture soma_sub8 of soma_sub8 is
	-- <COMPLETAR>
begin

    -- <COMPLETAR>

end architecture;