--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

--------------------------------------
-- Entidade
--------------------------------------
entity soma_sub is
	port (-- <COMPLETAR>
	     );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture soma_sub of soma_sub is
	-- <COMPLETAR>
begin

    -- <COMPLETAR>
	
end architecture;