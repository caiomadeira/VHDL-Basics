--------------------------------------
-- Biblioteca
--------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--------------------------------------
-- Entidade
--------------------------------------
entity top is
	port (-- <COMPLETAR>
	     );
end entity;

--------------------------------------
-- Arquitetura
--------------------------------------
architecture top of top is
	-- <COMPLETAR>
begin

	-- <COMPLETAR>

end architecture;